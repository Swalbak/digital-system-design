library verilog;
use verilog.vl_types.all;
entity CH2_F_SEP_TB is
end CH2_F_SEP_TB;
