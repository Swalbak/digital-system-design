library verilog;
use verilog.vl_types.all;
entity CH2_4COMPARE_TB is
end CH2_4COMPARE_TB;
