library verilog;
use verilog.vl_types.all;
entity COUNT_8BIT_TB is
end COUNT_8BIT_TB;
