library verilog;
use verilog.vl_types.all;
entity ch2_18DEMUX_TB is
end ch2_18DEMUX_TB;
