library verilog;
use verilog.vl_types.all;
entity CH2_SYNC_3CNT2_TB is
end CH2_SYNC_3CNT2_TB;
