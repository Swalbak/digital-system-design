library verilog;
use verilog.vl_types.all;
entity CH2_BCDCONVERTER_TB is
end CH2_BCDCONVERTER_TB;
