library verilog;
use verilog.vl_types.all;
entity CH2_4PISO_TB is
end CH2_4PISO_TB;
