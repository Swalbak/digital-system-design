library verilog;
use verilog.vl_types.all;
entity CH2_83ENCODER_TB is
end CH2_83ENCODER_TB;
