library verilog;
use verilog.vl_types.all;
entity CH2_2MUX_TB is
end CH2_2MUX_TB;
